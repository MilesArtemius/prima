�� sr classes.graph.Graph        L arkst Ljava/util/LinkedList;L nodest Ljava/util/HashMap;xpsr java.util.LinkedList)S]J`�"  xpw   sr classes.graph.Ark        Z hiddenD weightL endt Lclasses/graph/Node;L startq ~ xp@      sr classes.graph.Node        Z hiddenL arksq ~ L namet Ljava/lang/String;L positiont Ljava/awt/geom/Point2D;xpsq ~ w   q ~ sq ~ @      sq ~ 	sq ~ w   q ~ sq ~ @       sq ~ 	sq ~ w   q ~ sq ~ @      q ~ sq ~ 	sq ~ w   q ~ q ~ xt Asr java.awt.geom.Point2D$DoubleU[��	�_ D xD yxp@i      @y      xt Dsq ~ @@     @Y      q ~ xt Csq ~ @@     @��     q ~ xt Bsq ~ @�      @y      q ~ q ~ q ~ q ~ xsr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      q ~ q ~ q ~ q ~ q ~ q ~ q ~ q ~ x